*555 MCE
*Sngl Timer (Macromodel) pkg:DIP8 1,2,3,4,5,6,7,8
*Connections:
*              Gnd 
*              |  Trig
*              |  |  Out
*              |  |  |  Reset
*              |  |  |  |  Ctrl
*              |  |  |  |  |  Thresh
*              |  |  |  |  |  |  Dischg
*              |  |  |  |  |  |  |  Vcc
*              |  |  |  |  |  |  |  |
.SUBCKT 555    1  2  3  4  5  6  7  8 
EREF 15 1 8 1 .5
GSOURCE 8 3 8 26 12.5E-3
GSINK 3 1 26 1 67E-3
VD1 8 27 DC .8
VD2 28 1 DC .85
VREF 30 1 DC 1.2
C1 29 1 700E-15
RREF2 30 1 100E3
RREF 15 1 100E3
ROUT 3 1 100K
R1 6 1 500E9
R2 2 1 500E9
R3 8 5 75E3
R4 5 9 75E3
R5 9 1 75E3
R6 10 11 1E3
R7 13 14 1E3
R8 8 12 150E3
R9 4 8 500E9
R10 20 19 1E3
R11 16 17 1E3
R12 8 18 150E3
R13 8 21 150E3
R14 22 23 1E3
R15 8 26 150E3
R16 24 25 1E3
R19 7 1 500E9
R20 29 26 1E6
D1 1 11 DMOD
D2 12 11 DMOD
D3 12 14 DMOD
D4 1 14 DMOD
D5 18 17 DMOD
D6 1 17 DMOD
D7 18 19 DMOD
D8 1 19 DMOD
D9 21 14 DMOD
D10 21 25 DMOD
D11 1 23 DMOD
D12 18 23 DMOD
D13 26 25 DMOD
D14 1 25 DMOD1
D15 3 27 DMOD
D16 28 3 DMOD
E1 10 1 6 5 1000
E2 13 1 2 9 1000
E3 16 1 15 12 1000
E4 22 1 15 21 1000
E5 24 1 15 18 1000
E7 20 1 4 30 1000
M1 7 29 1 1 MOSMOD
.MODEL MOSMOD NMOS (LEVEL=1 KP=1 VTO=1 RD=5)
.MODEL DMOD D (RS=1E-6)
.MODEL DMOD1 D (RS=1E-6 IS=1E-9)
.ENDS 555
* Motorola IP=.5U IV=6M VB1(sat)=3 Rbb=6.1K Vob1=3.6: E, B1, B2
*Connections:
*              E
*              | B1
*              | | B2
*              | | |
.SUBCKT 2N2646 1 2 3
DE 1 4 EMITTER
VE 4 5 DC 0
HVE 6 0 VE 1K
RVE 0 6 1MEG
BBB 5 7 I=0.00028*V(5,7)+0.00575*V(5,7)*V(6)
CBB 5 7 35P
RB1 7 2 38.15 RMOD
RB2 3 5 2.518K RMOD 
.MODEL RMOD R TC1=.01
.MODEL EMITTER D (IS=21.3P N=1.8)
.ENDS 2N2646
------------------------------------------------------------
-- VHDL FPGAProject_Top
-- 2006 9 7 17 14 18
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2004 Altium Limited"
------------------------------------------------------------

------------------------------------------------------------
-- VHDL FPGAProject_Top
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity FPGAProject_Top Is
  attribute MacroCell : boolean;

End FPGAProject_Top;
------------------------------------------------------------

------------------------------------------------------------
architecture structure of FPGAProject_Top is


begin
end structure;
------------------------------------------------------------


.SUBCKT ETABLE 1 2 3 4
  E1 3 4 TABLE {V(1, 2)} = (2,3)(4,5)(6,7)(8,9)(10,11)(12,13)(14,12)(16,11)(18,10)(20,14)
.ENDS ETABLE














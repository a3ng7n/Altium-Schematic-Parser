*Unary Minus of Voltage
.SUBCKT UNARYV 1 2
BX 2 0 V=-(V(1))
.ENDS UNARYV
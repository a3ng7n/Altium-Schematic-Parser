*Vacuum Tube Triode (Audio freq.)
*Connections:
*             Plate
*             | Grid
*             | | Cathode
*             | | |
.SUBCKT 7199T 1 3 4
B1 2 4 I=((URAMP((V(2,4)/17)+V(3,4)))^1.5)/711
C1 3 4 2.3E-12
C2 3 1 2.0E-12
C3 1 4 0.3E-12
R1 3 5 5E+3
D1 1 2 DX
D2 4 2 DX2
D3 5 4 DX
.MODEL DX D(IS=1.0E-12 RS=1.0)
.MODEL DX2 D(IS=1.0E-9 RS=1.0)
.ENDS 7199T
